module pref

[heap]
pub struct Preferences {
pub mut:
	is_strict       bool
	suppress_output bool
}
