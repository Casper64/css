module datatypes

pub struct CalcSum {
}

// evaluate returns evaluates the sum and returns the value in pixels
pub fn (sum CalcSum) evaluate(em f64, rem f64, vh f64, vw f64) f64 {
	return 0.0
}
