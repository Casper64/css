module datatypes

pub struct CalcSum {
}

// evaluate returns evaluates the sum and returns the value in pixels
pub fn (sum CalcSum) evaluate(em f32, rem f32, vh f32, vw f32) f32 {
	return 0.0
}
